`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/07/19 20:55:09
// Design Name: 
// Module Name: knight_rider_test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module knight_rider_test(

    input clk,
    output [7:0] led_out
    );

    parameter LEDS_INIT = 10'b1100000000;
    parameter DIR_INIT = 1;

endmodule
